module top8227 (


);




endmodule