`include "param_file.sv"

module  (
    ports
);
    
endmodule