module programCH (
    input logic [7:0] ADH_in,
    input logic nrst, clk,
    input logic PCH_PCH,
    input logic ADH_PCH,
    input logic PCLC,
    input logic PCH_DB,
    input logic PCH_ADH,
    output logic [7:0] DB_out, ADH_out  //
);

endmodule